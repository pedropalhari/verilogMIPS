library verilog;
use verilog.vl_types.all;
entity cpu_TB is
end cpu_TB;
