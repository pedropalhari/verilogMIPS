library verilog;
use verilog.vl_types.all;
entity reg32bits_TB is
end reg32bits_TB;
