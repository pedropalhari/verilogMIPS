library verilog;
use verilog.vl_types.all;
entity registerfile_TB is
end registerfile_TB;
