library verilog;
use verilog.vl_types.all;
entity pc_TB is
end pc_TB;
