library verilog;
use verilog.vl_types.all;
entity extend_TB is
end extend_TB;
